

module im_4k_test();
reg [31:0]addr;
wire [31:0] dout;
im_4k dd(addr,dout);
initial 
begin
#0 addr =32'b00000000000000000000000000000001+32'o0000_3000;
#10 addr=32'b00000000000000000000000000000010+32'o0000_3000;
#30 addr=32'b00000000000000000000000000000011+32'o0000_3000;
end
endmodule