library verilog;
use verilog.vl_types.all;
entity test_Risc_16_bit is
end test_Risc_16_bit;
