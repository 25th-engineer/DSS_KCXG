library verilog;
use verilog.vl_types.all;
entity mux_tb is
end mux_tb;
