library verilog;
use verilog.vl_types.all;
entity tb_mips16 is
end tb_mips16;
