library verilog;
use verilog.vl_types.all;
entity Risc_16_bit is
    port(
        clk             : in     vl_logic
    );
end Risc_16_bit;
