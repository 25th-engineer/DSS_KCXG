`include "npc.v"
`include "pc.v"
`include "regfile.v"
`include "ALU.v"
`include "signext.v"
`include "dm_4k.v"
`include "mux.v"
`include "im_4k.v"
`include "trancode.v"
module datapath(pc,npc,busA,busB,result,inscode,clk,rst,op,func,regdst,ALUsrc,memtoreg,regwr,memwr,branch,jump,ALUop,extop,extout,dmout,mux_result,mux2_data,imm16,rs,rt,rd,Target,zero);
input clk,rst ;
input [31:0]pc,inscode;
input regdst,ALUsrc,memtoreg,regwr,memwr,branch,jump,extop;
input [2:0]ALUop;
input [31:0]npc;
input zero;
output wire [5:0]op,func;
input [31:0] busA,busB,result;//,inscode;
wire [31:0]imm32;
input [31:0] extout,dmout,mux_result,mux2_data;
input [15:0] imm16;
input [4:0]rs,rt,rd;
input [25:0] Target;
/*module ALU(
input [2:0] ALUctr,
input [32:0] rs, rt,
output zero,
output reg [32:0] ALUout
);  */
ALU alu(ALUop,busA,mux_result,zero,result);
/*module PC(npc,clk,rst,pc);
input clk;
input rst;
input [31:0] npc;
output reg [31:0] pc;*/
pc per_pc(npc,clk,rst,pc);
/*
module npc(zero,branch,Imm16,pc,npcTarget,jump);
input zero ;
input branch ;  
input [31:0] pc ;
input [15:0] Imm16;
output [31:0] npc;
*/
npc next_pc (zero,branch,imm16,pc,npc,Target,jump);

/*module im_4k(
input [31:0] addr,
output reg [31:0] dout);*/
im_4k instrution( pc,inscode);
/*module trancode (inscode,op,rs,rt,rd,Target,imm16);
*/
trancode code(inscode,op,rs,rt,rd,Target,imm16,func);

/*module mux #(parameter WIDTH = 32) 
(input [WIDTH-1:0] d0, d1,	
	input s,		
	output [WIDTH-1:0] y);	
*/
mux mux2(busB,extout,ALUsrc,mux_result);

/*module dm_4k (
input [11:2]addr,
input [31:0] din,
input we,
input clk,
output [31:0] dout
);*/
dm_4k datamem(result,busB,memwr,clk,dmout);
mux mux2_2(result,dmout,memtoreg,mux2_data);

/*module regfile(
input clk,
input [4:0] rd,rs,rt,
input [31:0]busw,
output [31:0]busA,busB,
input regwr,regdst
);*/

regfile registerfile(clk,rd,rs,rt,mux2_data,busA,busB,regwr,regdst);

/*module signext #(parameter WIDTH=16)(
input [WIDTH-1:0]imm16,
input extop,
output reg[31:0]imm32);*/
signext ext(imm16,extop,extout);
signext ex(imm16,1,imm32);

endmodule 
